module hello;
    initial
        $display("Hello!");
endmodule
