module hello_world;
  initial
    $display("Hello World !");
endmodule
