module main;
    hello my_hello();
    hello my_hello2();

    initial
    begin
        $display("test");
    end
endmodule
